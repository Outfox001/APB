// ---------------------------------------------------------------------------------------------------------------------
// Module name: afvip_intrr_pkg
// HDL        : System Verilog
// Author     : Paulovici Vlad-Marian
// Description: Package for signal interrupt
// Date       : 28 August, 2023
// ---------------------------------------------------------------------------------------------------------------------
package afvip_intrr_pkg;

  import uvm_pkg::*;

  `include "uvm_macros.svh"
  `include "afvip_intrr_item.svh"
  `include "afvip_intrr_monitor.svh"
  `include "afvip_intrr_agent.svh"
  `include "afvip_intrr_coverage.svh"

endpackage