// ------------------------------------------------------------------------------------------------------------------------------------------------------------------------
// Module name: afvip_test_pkg
// HDL        : UVM
// Author     : Paulovici Vlad-Marian
// Description: Package for the library of tests and virtual sequence
// Date       : 28 August, 2023
// -----------------------------------------------------------------------------------------------------------------------------------------------------------------------------


package afvip_test_pkg;

  import uvm_pkg::*;
  import afvip_apb_pkg::*;
  import afvip_reset_pkg::*;
  import afvip_intrr_pkg::*;
  import afvip_env_pkg::*;

  `include "uvm_macros.svh"
  `include "afvip_test_lib.svh"
   
endpackage